module part3(
  input A[3:0],B[3:0],OPCODE[2:0],
  output Y[3:0],N,Z,C,V
  );
endmodule
